module datapath(
	//input logic[15:0] S,
);



endmodule