module reg_file
(input logic [2:0] DR, SR2, SR1
 input logic LD_REG, Clk
);

R1

endmodule
