module register_unit(
)



endmodule